

/*

Converts a four-bit binary number V = v3v2v1v0 into a two-digit decimal equivalent D = d1d0. 
For example, if the input (V = 1111), then we would get 15 as the output in the 7-segment display. 
Use a comparator to check when the value of V is greater than 9, 
and use the output of this comparator in the control of the 7-segment displays. 


*/ 


